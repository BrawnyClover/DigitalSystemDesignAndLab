module temp(
inp1, out1
);

input [6:0] inp1;
output wire [6:0] out1;

assign out1 = inp1;

endmodule
